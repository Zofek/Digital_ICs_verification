`timescale 1ns/1ps

package mult_pkg;
	
    import uvm_pkg::*;
`include "uvm_macros.svh"

//------------------------------------------------------------------------------
// package typedefs
//------------------------------------------------------------------------------

	typedef enum bit[2:0] {
		RST_OP        = 3'b000,
		CORR_INPUT    = 3'b001,
		INCORRECT_A   = 3'b010,
		INCORRECT_B   = 3'b011,
		INCORRECT_A_B = 3'b100
	} operation_t;
	
    // terminal print colors
    typedef enum {
        COLOR_BOLD_BLACK_ON_GREEN,
        COLOR_BOLD_BLACK_ON_RED,
        COLOR_BOLD_BLACK_ON_YELLOW,
        COLOR_BOLD_BLUE_ON_WHITE,
        COLOR_BLUE_ON_WHITE,
        COLOR_DEFAULT
    } print_color;

//    // WRITE COMMAND data packet
//    typedef struct packed 
//    {	
//		shortint 	arg_a;
//	    shortint 	arg_b;
//		bit 		arg_a_parity;
//		bit 		arg_b_parity;
//	    operation_t op;
//    } command_s;
	
	// WRITE RESULT data packet
//	typedef struct packed 
//	{
//		bit 	arg_parity_error;
//		int 	result;
//		bit 	result_parity; 					
//
//	} result_s;

//------------------------------------------------------------------------------
// package functions
//------------------------------------------------------------------------------

    // used to modify the color of the text printed on the terminal

    function void set_print_color ( print_color c );
        string ctl;
        case(c)
            COLOR_BOLD_BLACK_ON_GREEN : ctl  = "\033\[1;30m\033\[102m";
            COLOR_BOLD_BLACK_ON_RED : ctl    = "\033\[1;30m\033\[101m";
            COLOR_BOLD_BLACK_ON_YELLOW : ctl = "\033\[1;30m\033\[103m";
            COLOR_BOLD_BLUE_ON_WHITE : ctl   = "\033\[1;34m\033\[107m";
            COLOR_BLUE_ON_WHITE : ctl        = "\033\[0;34m\033\[107m";
            COLOR_DEFAULT : ctl              = "\033\[0m\n";
            default : begin
                $error("set_print_color: bad argument");
                ctl                          = "";
            end
        endcase
        $write(ctl);
    endfunction

//------------------------------------------------------------------------------
// testbench classes
//------------------------------------------------------------------------------	
	`include "random_command_transaction.svh"
	`include "minmax_command_transaction.svh"
	`include "result_transaction.svh"	
	`include "coverage.svh"
	`include "tpgen.svh"
	`include "scoreboard.svh"
	`include "driver.svh"
	`include "command_monitor.svh"
	`include "result_monitor.svh"
	`include "env.svh"
//------------------------------------------------------------------------------
// test classes
//------------------------------------------------------------------------------
	`include "random_test.svh"
	`include "minmax_test.svh"

endpackage : mult_pkg
